module main

// Coord holds a position within 2d space
struct Coord {
	x int
	y int
}