module main

// Coord holds a position within 2d space
struct Coord {
mut:
	x int
	y int
}