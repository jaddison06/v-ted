module main

struct Coord {
	x int
	y int
}