module main

fn main() {
	mut app := &App{}
	app.init("../main.v.bak")
	app.start()?
}

// todo:
//   -> menu impl
//   -> allow side-by-side menu options as well as vertical
//   -> scrolling
//   -> cursor move
//   -> typing, backspace, etc (elegant impl PLEASE)
//   -> ctrl+q to quit, ctrl+alt+q to force
//        -> get rid of esc to quit - instead we can use that to exit menus,
//           multiple cursors, other contextual stuff
//   -> save file (& warning menu on close w/o save)
//   -> ctrl+(shift|alt)+s to save as new file
//   -> start empty, ctrl+o to open file
//   -> multiple files in different tabs
//        -> scrollable on overflow
//        -> drag/drop to reorder, divider becomes bold at insert location
//   -> ctrl+n for new file, when saved it goes to save as
//   -> command line arg parser
//   -> scroll bar
//   -> highlighting
//   -> copy/paste w/ v clipboard lib
//   -> syntax highlighting w/ textmate
//   -> workspace file browser
//   -> ctrl+f to find in file, ctrl+(shift|alt)+f to find in workspace
//   -> ctrl+(shift|alt)+o to open new workspace (closes the current one)
//   -> find yaml lib? or write one it can't be that hard...
//   -> <home>/.vcoder/config.yaml
//   -> platform-independent settings module - can find "home" dir
//   -> settings menu
//        -> text tab format (tabs/spaces)
//             -> impl rendering tabs as spaces, but saving as tabs
//             -> vs code will shit itself - enforce spaces? -> space count is configurable
//        -> pre-written commands
//   -> ctrl+r to run pre-written command, ctrl+(shift|alt)+r to run arbitrary (output where?)
//   -> editing extras
//        -> ctrl+backspace to delete word
//        -> shift+cursor move to highlight (works w/ end, home, up, down, etc)
//        -> multiple cursors?
//             -> alt-click to add new
//             -> configurable blink speed
//             -> hide actual term cursor, instead highlight & blank characters